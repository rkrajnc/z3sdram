module cs8900a_8bit (
	clk,
	reset,
	en,
	nIOR,
	nIOW,
	addr
	
);

input clk;
input reset;
input en;
input nIOR;
input nIOW;
input [3:0] addr;


always @(posedge clk) begin
	
end

endmodule